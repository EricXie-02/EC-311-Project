`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/19/2022 07:57:44 PM
// Design Name: 
// Module Name: SSD_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SSD_test(
    input [1:0] state
    );
    reg SSD_A,SSD_B,SSD_C,SSD_D,SSD_E;
endmodule
